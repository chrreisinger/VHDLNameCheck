package alutb is
end alutb;

package body alutb is
  --constant foo_bar : integer;
  --variable x       : real;
  --type     myInt is range 0 to 10;

  function foodf (
    constant foo : integer)
    return integer is
  begin  -- foo_df
  end foodf;

end alutb;
