package alutb is
end alutb;

package body alutb is
  --constant foo_bar : integer;
  --variable x       : real;
  --type     myInt is range 0 to 10;

  function foodf (
    constant foo : integer)
    return integer is
  begin  -- foo_df
    --CQDelay := SelectDelay((1 => (clk_ipd'last_event, tpd_clk_dataout_posedge, true)));
    --TODO Write(L, String'(" # Warning, "));
    --TODO l := new string'("");
    --TODO  Write (StrPtr5, STRING'( "(" ) );
    --return string'("?");
    report packagename'xeft severity note;
    x := 'x';
  end foodf;

end alutb;
